* This file contains all the subcircuits to be used in SRAM256.cir

***** long channel VTP = -0.9, VTN = 0.8 *****
*.include modelcard/1um.pm
*.param supply = 5
*.param ll = 1u

****** 50nm models***


.include 50nm-2.pm
.param supply =1

.param lambda=25nm
.param ll='2*lambda'

****** 16nm low power models***
*.include ./modelcard/PTM_LP/16nm.pm
*.param supply =0.9
*.param ll=16nm

****** 16nm high peformance models***
*.include ./modelcard/PTM_HP/16nm.pm
*.param supply =0.7
*.param ll=16nm


.subckt wire iot iof len=10 wid=10
*was rr=0.8 cc=200e-15
.param rr=0.4
.param cc = '100e-15'
rt iot iof 'rr*len*50/(wid)'
cf iof  0  'cc*len*wid*50/1e6'
.ends

.subckt wire_dual lt rt lf rf len=10 wid=10
Xt lt rt wire len='len' wid='wid'
Xf lf rf wire len='len' wid='wid'
.ends



.subckt nn d g s  ww=100
mnfet d g s 0 nmos L=ll w='ww*ll'
.ends

.subckt pp d g s   ww=100
mpfet d g s vdd pmos L=ll w='ww*ll'
.ends


.subckt inv out inn size=30 beta=2
XPP out inn vdd pp ww='size*beta/(beta+1)'
XNN out inn gnd nn ww='size/(beta+1)'
.ends

.subckt nnd2 out in1 in0 size=30 beta=2
Xap0 out in0 vdd pp ww='beta*size/(beta+2)'
Xap1 out in1 vdd pp ww='beta*size/(beta+2)'
Xan0 out in0 nng nn ww='2*size/(beta+2)'
Xan1 nng in1 0   nn ww='2*size/(beta+2)'
.ends nnd2

.subckt nor2 out in1 in0 size=30 beta=2
Xap0 ppi in0 vdd pp ww='2*beta*size/(2*beta+1)'
Xap1 out in1 ppi pp ww='2*beta*size/(2*beta+1)'
Xan0 out in0 0 nn ww='1*size/(2*beta+1)'
Xan1 out in1 0   nn ww='1*size/(2*beta+1)'
.ends nor2

.subckt latch out inn clk clb size=25 beta=2
Xn inn clk qin nn ww='5'
Xp inn clb qin pp ww='10'
Xfb qin ggg    inv size=10 beta=1
Xi ggg qin     inv size='size'
Xo out ggg     inv size='3*size'
.ends latch

.subckt flop qqq ddd clk
Xinve clb clk inv
Xflip int ddd clb clk latch
Xflop qqq int clk clb latch
.ends flop

.subckt reg8 ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0 in7 in6 in5 in4 in3 in2 in1 in0 clk
x7 ot7 in7 clk flop
x6 ot6 in6 clk flop
x5 ot5 in5 clk flop
x4 ot4 in4 clk flop
x3 ot3 in3 clk flop
x2 ot2 in2 clk flop
x1 ot1 in1 clk flop
x0 ot0 in0 clk flop
.ends reg8


* This buffers the output of a pulse source to give realistic edges
* It is defined to give a number of pulses, then stop
.subckt dat1 out period=1ns start=1ns sz=50 total=5 duty=3
V0 j0  0  PULSE('supply' 0 'start' 10p 10p 'duty*period' 'total*period')
x7 out j0 inv size='sz'
.ends dat1

*generates different data stream on all eight channels, buffered output
.subckt dat8 o7 o6 o5 o4 o3 o2 o1 o0 per=1ns start=1ns size=50
V0 j0  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' 'per')
V1 j1  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '2*per')
V2 j2  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '3*per')
V3 j3  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '4*per')
V4 j4  0  PULSE('supply' 0 'start' 10p 10p '0.5*per-10ps' '1*per')
V5 j5  0  PULSE('supply' 0 'start' 10p 10p '1*per-10ps' '2*per')
V6 j6  0  PULSE('supply' 0 'start' 10p 10p '1.5*per-10ps' '3*per')
V7 j7  0  PULSE('supply' 0 'start' 10p 10p '2*per-10ps' '4*per')
xb o7 o6 o5 o4 o3 o2 o1 o0 j7 j6 j5 j4 j3 j2 j1 j0 buf8 sz='size'
.ends dat8

.subckt buf8 ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0 in7 in6 in5 in4 in3 in2 in1 in0 sz=100
x7 ot7 in7 inv size='sz'
x6 ot6 in6 inv size='sz'
x5 ot5 in5 inv size='sz'
x4 ot4 in4 inv size='sz'
x3 ot3 in3 inv size='sz'
x2 ot2 in2 inv size='sz'
x1 ot1 in1 inv size='sz'
x0 ot0 in0 inv size='sz'
.ends buf8


.subckt nnd3 out in2 in1 in0 size=20 beta=2
Xp0 out in0 vdd pp ww='beta*size/(beta+3)'
Xp1 out in1 vdd pp ww='beta*size/(beta+3)'
Xp2 out in2 vdd pp ww='beta*size/(beta+3)'
Xn0 out in0 nn0 nn ww='3*size/(beta+3)'
Xn1 nn0 in1 nn1 nn ww='3*size/(beta+3)'
Xn2 nn1 in2 gnd nn ww='3*size/(beta+3)'
.ends

.subckt senseAmp ot1 ot0 in1 in0 eva size=40
Xn0 ot0 in0 ot1 eva nnd3 size ='size'
Xn1 ot1 in1 ot0 eva nnd3 size ='size'
.ends senseAmp


* model for a single bit or memory
.subckt mem1 it if ac
xpst it ac tt  nn ww=5
xpsf if ac ff  nn ww=5
Xpif tt ff vdd pp ww=5
xpit ff tt vdd pp ww=5
Xnit tt ff gnd nn ww=5
xnif ff tt gnd nn ww=5
.ends mem1




* The critical path logic for the decoder is placed in here
* it uses just a single bit
* It is only necessary to model the worst case path through the logic
* Wire models are not necessary here, but be aware that wires might be
*significant in a real design
.subckt decodeModel choose Din clk sz=100
Xn0 dinf Din inv

Xn1 i1 dinf vdd nnd2
Xn2 ded1 dinf gnd nnd2

Xn3 i2 i1 gnd nor2
Xn4 ded2 i1 vdd nor2

Xn5 i3 i2 vdd nnd2
Xn6 ded3 i2 gnd nnd2

Xn7 i4 i3 inv

Xn8 i5 i3 clk nnd2

Xn9 choose i5 inv
.ends decodeModel


*Place the circuit to write the bit lines here
* btt and bff are the bit lines that must be reset when clk=LO
* dii is the value to be written
* rwt chooses either to read or write
* both dii and rwt must be timed through flop
.subckt write1 btt bff dii rwt clk sz=100
Xiclk clkf clk inv

Xnor2 wrt rwt clkf nor2

Xtn1 i1 wrt gnd nn
Xtn2 btt dii i1 nn
xtp3 vdd wrt btt pp

Xidi diif dii inv

Xtn4 bff diif i1 nn
Xtn5 vdd wrt bff pp
.ends write1


*Place the circuit to read the bit lines here
* btt and bff are the bit lines that must be reset when clk=LO
* out is the value read, it must be clocked into flop
* rwt chooses either to read or write
*
** you can use the subck 'senseAmp' if desired
.subckt read1 btt bff out rwt clk
Xn0 rd rwt clk nnd2
Xn1 rdf rd inv

Xn2 reset btt set rdf nnd3 size =40
Xn3 set bff reset rdf nnd3 size =40

Xn4 resetf reset inv

Xn5 setf set inv
Xn6 setff setf inv

Xn7 vdd setff i1 pp
Xn8 i1 resetf gnd nn

Xn9 out i1 inv
Xn10 i1 out inv
.ends read1



